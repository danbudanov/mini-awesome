/**
* @file ADS1672_EVM_tb.sv
* @author Daniil Budanov
* @brief Testbench for the ADS1672-EVM ADC
*/

module ADS1672_EVM_tb;
endmodule
